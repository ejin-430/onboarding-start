`default_nettype none
`timescale 1ns / 1ps

/* This testbench just instantiates the module and makes some convenient wires
   that can be driven / tested by the cocotb test.py.
*/
module tb ();

  // Dump the signals to a VCD file. You can view it with gtkwave or surfer.
  initial begin
    $dumpfile("tb.vcd");
    $dumpvars(0, tb);
    #1;
  end

  // Wire up the inputs and outputs:
  reg clk;
  reg rst_n;
  reg ena;
  reg [7:0] ui_in;
  reg [7:0] uio_in;
  wire [7:0] uo_out;
  wire pwm_out;
  assign pwm_out = uo_out[0];
  wire [7:0] uio_out;
  wire [7:0] uio_oe;
  
  // Give reg inputs a known value at time 0 (avoids Xs in gate-level sim)
  initial begin
    clk    = 1'b0;
    rst_n  = 1'b1;
    ena    = 1'b0;
    uio_in = 8'h00;

    // SPI idle (Mode 0): nCS=1, COPI=0, SCLK=0
    // ui_in[2]=nCS, ui_in[1]=COPI, ui_in[0]=SCLK  => 0b00000100
    ui_in  = 8'h04;
  end

`ifdef GL_TEST
  wire VPWR = 1'b1;
  wire VGND = 1'b0;
`endif

  // Replace tt_um_example with your module name:
  tt_um_uwasic_onboarding_eva_jin user_project (

      // Include power ports for the Gate Level test:
`ifdef GL_TEST
      .VPWR(VPWR),
      .VGND(VGND),
`endif

      .ui_in  (ui_in),    // Dedicated inputs
      .uo_out (uo_out),   // Dedicated outputs
      .uio_in (uio_in),   // IOs: Input path
      .uio_out(uio_out),  // IOs: Output path
      .uio_oe (uio_oe),   // IOs: Enable path (active high: 0=input, 1=output)
      .ena    (ena),      // enable - goes high when design is selected
      .clk    (clk),      // clock
      .rst_n  (rst_n)     // not reset
  );

endmodule
